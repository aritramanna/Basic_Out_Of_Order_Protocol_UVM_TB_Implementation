package axi_uvm_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "transaction.sv"
`include "sequence.sv"
`include "wr_rd_sequence_random_id.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "env.sv"
`include "test.sv"

endpackage