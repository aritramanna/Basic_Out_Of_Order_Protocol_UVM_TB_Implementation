
`include "ooo_pkg.sv"
`include "interface.sv"
`include "tb.sv"
